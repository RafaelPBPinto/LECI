library ieee;
use ieee.std_logic_1164.all;

entity Dec2_4ENDemo is
	port (SW  : in std_logic_vector(2 downto 0);
			LedG: out std_logic_vector(3 downto 0));
end Dec2_4ENDemo;

architecture Shell of Dec2_4EnDemo is
begin
	system_core : work entity.Dec2_4En(BehavEquations)
		port map(enable <= SW(2);
					inputs <= SW;
					outputs => LedG(3 downto 0));
end Dec2_4EnDemo;	