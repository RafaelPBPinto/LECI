library ieee;
use ieee.std_logic_1164.all;

entity latch1 is 
	port (enable : in std_logic;
			d      : in std_logic;
			q      : out std_logic);
end latch1;

architecture v1 of latch1 is

begin 
	process(enable)
	begin
		if(enable = '1') then
			q <= d;
		end if;
	end process;
end v1;